*sumator.spi
* Netlista sumatora
.subckt SUMATOR A B C SUM CARRY VDD VSS


********************Blok CARRY
*Tablica PMOS
M1 s1 A VDD VDD PCH L=0.065u W=0.94u M=1
M2 s1 B VDD VDD PCH L=0.065u W=0.94u M=1
M3 s2 B s1 VDD PCH L=0.065u W=0.94u M=1
M4 Ca C s1 VDD PCH L=0.065u W=0.94u M=1
M5 Ca A s2 VDD PCH L=0.065u W=0.94u M=1

*Tablica NMOS
M6 Ca C s3 VSS NCH L=65n W=200n M=1
M7 Ca A s4 VSS NCH L=65n W=200n M=1
M8 s3 A VSS VSS NCH L=65n W=200n M=1
M9 s3 B VSS VSS NCH L=65n W=200n M=1
M10 s4 B VSS VSS NCH L=65n W=200n M=1

*INV
M11 CARRY Ca VDD VDD PCH L=0.065u W=0.94u M=1
M12 CARRY Ca VSS VSS NCH L=65n W=200n M=1

********************BLOK SUM
*Tablica PMOS
M13 s5 A VDD VDD PCH L=0.065u W=0.94u M=1
M14 s5 B VDD VDD PCH L=0.065u W=0.94u M=1
M15 s5 C VDD VDD PCH L=0.065u W=0.94u M=1
M16 s6 A s5 VDD PCH L=0.065u W=0.94u M=1
M17 s7 B s6 VDD PCH L=0.065u W=0.94u M=1
M18 S C s7 VDD PCH L=0.065u W=0.94u M=1
M19 S Ca s5 VDD PCH L=0.065u W=0.94u M=1

*Tablica NMOS

M20 s8 A VSS VSS NCH L=65n W=200n M=1
M21 s8 B VSS VSS NCH L=65n W=200n M=1
M22 s8 C VSS VSS NCH L=65n W=200n M=1
M23 s9 B VSS VSS NCH L=65n W=200n M=1
M24 s10 A s9 VSS NCH L=65n W=200n M=1
M25 S C s10 VSS NCH L=65n W=200n M=1
M26 S Ca s8 VSS NCH L=65n W=200n M=1


*INV
M27 SUM S VDD VDD PCH L=0.065u W=0.94u M=1
M28 SUM S VSS VSS NCH L=65n W=200n M=1

.ends