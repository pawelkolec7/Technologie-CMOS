.INCLUDE sumator.spi

xSUMATOR1 VDD VSS C0 SUM0 CARRY0 VDD VSS SUMATOR
xSUMATOR2 VDD VSS CARRY0 SUM1 CARRY1 VDD VSS SUMATOR
xSUMATOR3 VDD VSS CARRY1 SUM2 CARRY2 VDD VSS SUMATOR
xSUMATOR4 VDD VSS CARRY2 SUM3 CARRY3 VDD VSS SUMATOR
* Supply DC voltage

VDD VDD VSS DC 1.2
VSS VSS 0 0

* Source(LOW HIGH DELAY RISE FALL WIDTH PERIOD)

VC0 C0 VSS PULSE (0.0 1.2 0.0 0.01n 0.01n 1n 2n)

* Load

.end